module project6(

   );
endmodule