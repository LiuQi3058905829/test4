module D(

   );
endmodule