module D1(

   );
endmodule