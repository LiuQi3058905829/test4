module AyB(

   );
endmodule