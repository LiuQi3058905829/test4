module gate74LS74(

   );
endmodule